** Profile: "SCHEMATIC1-sim"  [ D:\facultate\an_3\sem_1\proiect apd_proiect cef\P1_2024_431A_Sava_Rares_PACT_N10_OrCAD\Schematics\schema_electronica-pspicefiles\schematic1\sim.sim ] 

** Creating circuit file "sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../lib_modelespice/lib_modelepspice_anexa_1/modele_a1_lib/bc807-25.lib" 
.LIB "../../../lib_modelespice/lib_modelepspice_anexa_1/modele_a1_lib/bc817-25.lib" 
.LIB "../../../lib_modelespice/lib_modelepspice_anexa_1/modele_a1_lib/bc846b.lib" 
* From [PSPICE NETLIST] section of C:\Users\rares\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.AC DEC 10 1 1Meg
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
